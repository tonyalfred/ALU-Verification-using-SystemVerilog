`include "alu_if.sv"

package env_pkg; 
	`include "packet.svh"
	`include "scoreboard.svh"
	`include "monitor.svh"
	`include "driver.svh"
	`include "stimulus_gen.svh"
endpackage 